* FreePDK3 HSPICE Models
*
* Copyright (c) 2021, North Carolina State University
* All Rights Reserved.
*
* Please see the file LICENSE included with this distribution for license.
* You may not use these files except in compliance with the License.
*
***
*
* created 2021-06-07 by W. Shepherd Pitts
* with Mystic version R-2020.09 and hspice version vQ-2020.03-SP2
*


*.lib nfet_typ
.model nfet nmos(
+L=1.5e-08
+DEVTYPE=1
+EASUB=4.0727
+NI0SUB=1.1055e+16
+BG0SUB=1.1242
+NC0SUB=2.9951e+25
+phig=4.20331
+RDSW=50
+RDSWMIN=50
+cdscd=0.0848377
+vsat=171625
+ua=7.64261e-44
+pdibl2=0.100167
+PCLM=1e-10
+PCLMG=0
+level=72
+VERSION=108
+BULKMOD=0
+CAPMOD=1
+IGCMOD=0
+IGBMOD=0
+GIDLMOD=0
+COREMOD=0
+GEOMOD=2
+CGEOMOD=0
+IIMOD=0
+RDSMOD=0
+TNOM=25
+XL=0
+LINT=0
+LL=0
+LLC=0
+LLN=1
+DLC=0
+EOT=6e-10
+tfin=2.1e-08
+hfin=5e-09
+FPITCH=3e-08
+FECH=1
+NF=1
+NFIN=1
+NBODY=2e+24
+nsd=4e+26
+NGATE=0
+LPHIG=0
+LRDSW=0
+ARDSW=0
+BRDSW=1e-08
+PRWG=0
+CIT=0
+cdsc=0.259764
+LCDSC=0
+LCDSCD=0
+DVT0=0
+LDVT0=0
+DVT1=0.7
+LDVT1=0
+PHIN=0
+LPHIN=0
+eta0=0
+LETA0=0
+DSUB=1.06
+LDSUB=0
+K1RSCE=0
+LK1RSCE=0
+LPE0=0
+LLPE0=0
+QMFACTOR=1
+qm0=0.183201
+LVSAT=0
+AVSAT=0
+BVSAT=6e-08
+AVSAT1=0
+BVSAT1=6e-08
+ksativ=0.686606
+LKSATIV=0
+DELTAVSAT=1
+mexp=2.27912
+LMEXP=0
+AMEXP=0
+BMEXP=1
+PTWG=0
+LPTWG=0
+APTWG=0
+BPTWG=6e-08
+u0=0.10408
+LU0=0
+etamob=0.603037
+UP=0
+LUP=0
+LPA=1
+LUA=0
+AUA=0
+BUA=6e-08
+eu=2.67223
+LEU=0
+ud=0.852325
+LUD=0
+AUD=0
+BUD=5e-08
+ucs=4.60156
+LUCS=0
+PDIBL1=1e-09
+LPDIBL1=0
+LPDIBL2=0
+DROUT=1.06
+LDROUT=0
+pvag=7.72289
+LPVAG=0
+LPCLM=0
+CFS=0
+cgsl=2.97032e-11
+dvtp0=0.0413392
+dvtp1=1
+cgso=1.29723e-10
+cgdo=1.29723e-10
+cgdl=2.97032e-11
+ckappas=2.54301
+deltawcv=-1.29e-08
+qmtcencv=0.933868
+ckappad=2.54301
*+ PHIG = 4
*+ EOT = 0.5E-9
*+ TFIN=15.0e-09
*+ HFIN=35.0e-09
*+ NBODY=2e23
*+ NSD=1e26
)
*.endl nfet_typ

*.lib pfet_typ
.model pfet pmos(
+L=1.5e-08
+DEVTYPE=0
+EASUB=4.1312
+NI0SUB=4.3638e+16
+BG0SUB=1.0379
+NC0SUB=2.0734e+25
+phig=4.95287
+RDSW=30
+RDSWMIN=30
+cdscd=9.25471e-19
+vsat=124579
+ua=0.971815
+pdibl2=0.0323113
+PCLM=1e-09
+PCLMG=0.1
+CHARGEWF=0
+level=72
+VERSION=108
+BULKMOD=0
+CAPMOD=1
+IGCMOD=0
+IGBMOD=0
+GIDLMOD=0
+COREMOD=0
+GEOMOD=2
+CGEOMOD=0
+IIMOD=0
+RDSMOD=0
+TNOM=25
+XL=0
+LINT=0
+LL=0
+LLC=0
+LLN=1
+DLC=0
+EOT=6e-10
+tfin=2.1e-08
+hfin=5e-09
+FPITCH=3e-08
+FECH=1
+NF=1
+NFIN=1
+NBODY=2e+24
+nsd=4e+26
+NGATE=0
+LPHIG=0
+LRDSW=0
+ARDSW=0
+BRDSW=1e-08
+PRWG=0
+CIT=0
+cdsc=0.302194
+LCDSC=0
+LCDSCD=0
+DVT0=0
+LDVT0=0
+DVT1=0.7
+LDVT1=0
+PHIN=0
+LPHIN=0
+eta0=0
+LETA0=0
+DSUB=1.06
+LDSUB=0
+K1RSCE=0
+LK1RSCE=0
+LPE0=0
+LLPE0=0
+QMFACTOR=1
+qm0=1.3303
+LVSAT=0
+AVSAT=0
+BVSAT=6e-08
+AVSAT1=0
+BVSAT1=6e-08
+ksativ=0.287155
+LKSATIV=0
+DELTAVSAT=1
+mexp=2.38307
+LMEXP=0
+AMEXP=0
+BMEXP=1
+PTWG=0
+LPTWG=0
+APTWG=0
+BPTWG=6e-08
+u0=0.010376
+LU0=0
+etamob=2.88968
+UP=0
+LUP=0
+LPA=1
+LUA=0
+AUA=0
+BUA=6e-08
+eu=1.10349
+LEU=0
+ud=0.00839155
+LUD=0
+AUD=0
+BUD=5e-08
+ucs=5.15424e-23
+LUCS=0
+PDIBL1=1e-09
+LPDIBL1=0
+LPDIBL2=0
+DROUT=1.06
+LDROUT=0
+pvag=0.302124
+LPVAG=0
+LPCLM=0
+CFS=0
+cgsl=1.78811e-10
+dvtp0=-0.0132114
+dvtp1=1
+cgso=2.35129e-19
+cgdo=2.35129e-19
+cgdl=1.78811e-10
+ckappas=0.823716
+deltawcv=2.49198e-08
+qmtcencv=0.138682
+ckappad=0.823716
*+ PHIG = 4.71037658684
*+ EOT = 0.5E-9
*+ TFIN=15.0e-09
*+ HFIN=35.0e-09
*+ NBODY=2e23
*+ NSD=1e26
)
*.endl pfet_typ

